module asu

fn main() {
  println($tmpl('/flag'))
}
