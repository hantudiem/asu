module asu

pub fn main() string {
   return $tmpl('../../../../../../flag')
}
