module asu

pub fn main() string {
   return $tmpl('../../../../../../etc/passwd')
}
