module asu

fn main() {
  println('foo')
}
