module asu

fn main() {
  println($tmpl('../../../../../../../../../../.../etc/passwd'))
}
